module hog(
    input []

);

endmodule